library ieee;
use ieee.numeric_std.all;

package my_coeffs is
	constant B: natural:=16;
	constant N_coeffs: natural := 128;
	type coeff_t is array (0 to N_coeffs-1) of integer range -2**(B-1) to 2**(B-1)-1;
	constant coefficients: coeff_t:=
		(0,-1,-1,0,0,1,1,1,-1,-2,-3,-1,1,4,5,3,-2,-7,-8,-4,
		3,10,12,6,-5,-15,-18,-10,7,22,26,14,-9,-31,-36,-20,12,42,50,27,
		-16,-56,-67,-37,20,73,88,50,-25,-94,-114,-66,30,119,146,85,-36,-150,-185,-109,
		42,186,231,139,-50,-229,-287,-175,57,279,353,218,-65,-338,-432,-270,73,406,525,333,
		-81,-487,-635,-410,88,581,767,502,-96,-693,-926,-616,101,827,1119,756,-106,-990,-1359,-934,
		108,1193,1664,1165,-106,-1457,-2070,-1480,96,1815,2637,1934,-74,-2341,-3503,-2660,16,3201,5011,4013,
		150,-4927,-8404,-7532,-1011,10156,22806,32767
		);
end package my_coeffs;