library ieee;
use ieee.numeric_std.all;

package my_coeffs is
	constant B: natural:=16;
	constant N_coeffs: natural := 128;
	type coeff_t is array (0 to N_coeffs-1) of integer range -2**(B-1) to 2**(B-1)-1;
	constant coefficients: coeff_t:=
		(0,0,0,-1,-1,-1,0,2,2,2,1,-2,-4,-4,-3,1,5,8,7,2,
		-6,-11,-12,-7,3,14,20,17,4,-13,-26,-29,-17,6,29,42,35,10,-25,-53,
		-58,-35,10,56,81,69,20,-46,-98,-107,-65,16,100,144,123,37,-78,-168,-185,-113,
		24,165,241,206,66,-123,-273,-304,-188,33,261,385,332,111,-189,-426,-478,-301,42,399,
		596,520,181,-279,-649,-736,-472,50,598,907,802,293,-409,-981,-1129,-738,54,900,1392,1251,
		481,-608,-1517,-1780,-1196,46,1412,2247,2074,849,-964,-2553,-3102,-2181,-12,2543,4285,4191,1922,-1896,
		-5759,-7762,-6303,-755,8159,18463,27498,32767
		);
end package my_coeffs;