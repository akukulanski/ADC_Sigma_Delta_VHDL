package mytypes_pkg is
	type my_array_t is array (0 to 12) of natural; -- 12=2*N; N etapas
end package mytypes_pkg;