library ieee;
use ieee.numeric_std.all;

package my_coeffs is
	constant B: natural:=16;
	type coeff_t is array (TAPS-1 downto 0) of integer range -2**(B-1) to 2**(B-1)-1;
	constant coefficiets: coeff_t:=
		(0,0,0,0,1,1,1,0,-1,-2,-2,0,3,4,4,0,-4,-7,-6,-1,
		6,11,9,1,-10,-16,-14,-2,14,23,20,3,-19,-32,-28,-4,26,44,38,7,
		-34,-60,-51,-10,44,78,68,14,-57,-102,-89,-19,72,130,115,26,-90,-164,-146,-35,
		111,205,184,47,-135,-254,-229,-61,163,311,284,79,-196,-380,-350,-102,233,460,428,130,
		-277,-555,-521,-165,327,667,633,209,-385,-802,-769,-264,453,964,936,333,-534,-1164,-1145,-424,
		634,1416,1414,544,-760,-1747,-1775,-712,925,2203,2287,961,-1161,-2887,-3085,-1373,1529,4043,4519,2187,
		-2208,-6499,-7959,-4580,3821,15246,26139,32768
		);
end package my_coeffs;